package shared_pkg;
    typedef enum bit [1:0] {WR_ADDR, WR_DATA, RD_ADDR, RD_DATA } op_e;
endpackage
