package SPI_rd_only_sequence_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    import SPI_seq_item_pkg::*;
    import SPI_pkg::*;

    class SPI_rd_only_sequence extends uvm_sequence #(SPI_seq_item);
        `uvm_object_utils(SPI_rd_only_sequence)

        SPI_seq_item seq_item;

        function new(string name = "SPI_rd_only_sequence");
            super.new(name);
        endfunction

    task body();
        seq_item = SPI_seq_item::type_id::create("seq_item");
        //Read only
        repeat(5000) begin
            start_item(seq_item);
            //At the beginning of the operation, enable the read sequence and randomization
            if(counter_allcases == 0 && (seq_item.array_rand[0:2] inside {WR_ADDR, WR_DATA, RD_ADDR})
            || counter_read == 0 && (seq_item.array_rand[0:2] inside {RD_DATA})) begin
                seq_item.wr_only_constraint.constraint_mode(0);
                seq_item.rd_only_constraint.constraint_mode(1);
                seq_item.rd_wr_constraint.constraint_mode(0);            
                seq_item.array_rand.rand_mode(1);
            end
            else begin
                //Disable all constraints and randomization because we are already in an operation
                seq_item.wr_only_constraint.constraint_mode(0);
                seq_item.rd_only_constraint.constraint_mode(0);
                seq_item.rd_wr_constraint.constraint_mode(0);            
                seq_item.array_rand.rand_mode(0);
            end
            assert (seq_item.randomize());
            seq_item.update_counter_allcases;
            seq_item.update_counter_read;
            finish_item(seq_item);
        end

    endtask

endclass
endpackage