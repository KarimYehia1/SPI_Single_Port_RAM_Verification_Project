package shared_pkg;
int counter_allcases =0  ;
int counter_read=0;
 logic SS_n_prev=1;
endpackage