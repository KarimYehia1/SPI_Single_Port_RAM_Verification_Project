package SPI_SLAVE_shared_pkg;
typedef enum  {IDLE,CHK_CMD ,WRITE,READ_ADD , READ_DATA } current_st;
int counter_allcases =0  ;
int counter_read=0;
 logic SS_n_prev=1;
endpackage